-- Entitet: bitfeeder
-- Beskrivelse: Leverer to bit fra en fast defineret sekvens. Denne sekvens er et simuleret
-- SW kommunikationsflow (fra opstart til datatransmission). Her svarer bit1 til databit og bit0
-- til strobe. Dette skal simulere den kommunikationslinje systemet skal sidde på.

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity bit_feeder is
    Port (
        clk50mhz         : in  std_logic;
        reset       : in  std_logic;
        D     : out std_logic;
        S : out std_logic
    );
end entity;

architecture bit_feeder_arch of bit_feeder is

    -- Antallet af ROM elementer. Skal være stor nok til at kunne indeholde hele datapakken.
    constant ROM_SIZE : integer := 4000;

    -- Definerer ROM-typen som et array af 2-bit elementer
    type rom_type is array (0 to ROM_SIZE - 1) of std_logic_vector(1 downto 0);

    -- ROM-indhold: Forhåndsdefineret SW kommunikationsflow defineret som data og strobe
    
 constant rom : rom_type := (
	0 => "00", 1 => "00", 2 => "00", 3 => "00", 4 => "00", 5 => "00", 6 => "00", 7 => "00", 8 => "00", 9 => "00", 10 => "00", 11 => "00", 12 => "00", 13 => "00", 14 => "00", 15 => "00", 16 => "00", 17 => "00", 18 => "00", 19 => "00", 20 => "00", 21 => "00", 22 => "00", 23 => "00", 24 => "00", 25 => "00", 26 => "00", 27 => "00", 28 => "00", 29 => "00", 30 => "00", 31 => "00", 32 => "00", 33 => "00", 34 => "00", 35 => "00", 36 => "00", 37 => "00", 38 => "00", 39 => "00", 40 => "00", 41 => "00", 42 => "00", 43 => "00", 44 => "00", 45 => "00", 46 => "00", 47 => "00", 48 => "00", 49 => "00", 50 => "00", 51 => "00", 52 => "00", 53 => "00", 54 => "00", 55 => "00", 56 => "00", 57 => "00", 58 => "00", 59 => "00", 60 => "00", 61 => "00", 62 => "00", 63 => "00", 64 => "00", 65 => "00", 66 => "00", 67 => "00", 68 => "00", 69 => "00", 70 => "00", 71 => "00", 72 => "00", 73 => "00", 74 => "00", 75 => "00", 76 => "00", 77 => "00", 78 => "00", 79 => "00", 80 => "00", 81 => "00", 82 => "00", 83 => "00", 84 => "00", 85 => "00", 86 => "00", 87 => "00", 88 => "00", 89 => "00", 90 => "00", 91 => "00", 92 => "00", 93 => "00", 94 => "00", 95 => "00", 96 => "00", 97 => "00", 98 => "00", 99 => "00", 100 => "00", 101 => "00", 102 => "00", 103 => "00", 104 => "00", 105 => "00", 106 => "00", 107 => "00", 108 => "00", 109 => "00", 110 => "00", 111 => "00", 112 => "00", 113 => "00", 114 => "00", 115 => "00", 116 => "00", 117 => "00", 118 => "00", 119 => "00", 120 => "00", 121 => "00", 122 => "00", 123 => "00", 124 => "00", 125 => "00", 126 => "00", 127 => "00", 128 => "00", 129 => "00", 130 => "00", 131 => "00", 132 => "00", 133 => "00", 134 => "00", 135 => "00", 136 => "00", 137 => "00", 138 => "00", 139 => "00", 140 => "00", 141 => "00", 142 => "00", 143 => "00", 144 => "00", 145 => "00", 146 => "00", 147 => "00", 148 => "00", 149 => "00", 150 => "00", 151 => "00", 152 => "00", 153 => "00", 154 => "00", 155 => "00", 156 => "00", 157 => "00", 158 => "00", 159 => "00", 160 => "00", 161 => "00", 162 => "00", 163 => "00", 164 => "00", 165 => "00", 166 => "00", 167 => "00", 168 => "00", 169 => "00", 170 => "00", 171 => "00", 172 => "00", 173 => "00", 174 => "00", 175 => "00", 176 => "00", 177 => "00", 178 => "00", 179 => "00", 180 => "00", 181 => "00", 182 => "00", 183 => "00", 184 => "00", 185 => "00", 186 => "00", 187 => "00", 188 => "00", 189 => "00", 190 => "00", 191 => "00", 192 => "00", 193 => "00", 194 => "00", 195 => "00", 196 => "00", 197 => "00", 198 => "00", 199 => "00", 200 => "00", 201 => "00", 202 => "00", 203 => "00", 204 => "00", 205 => "00", 206 => "00", 207 => "00", 208 => "00", 209 => "00", 210 => "00", 211 => "00", 212 => "00", 213 => "00", 214 => "00", 215 => "00", 216 => "00", 217 => "00", 218 => "00", 219 => "00", 220 => "00", 221 => "00", 222 => "00", 223 => "00", 224 => "00", 225 => "00", 226 => "00", 227 => "00", 228 => "00", 229 => "00", 230 => "00", 231 => "00", 232 => "00", 233 => "00", 234 => "00", 235 => "00", 236 => "00", 237 => "00", 238 => "00", 239 => "00", 240 => "00", 241 => "00", 242 => "00", 243 => "00", 244 => "00", 245 => "00", 246 => "00", 247 => "00", 248 => "00", 249 => "00", 250 => "00", 251 => "00", 252 => "00", 253 => "00", 254 => "00", 255 => "00", 256 => "00", 257 => "00", 258 => "00", 259 => "00", 260 => "00", 261 => "00", 262 => "00", 263 => "00", 264 => "00", 265 => "00", 266 => "00", 267 => "00", 268 => "00", 269 => "00", 270 => "00", 271 => "00", 272 => "00", 273 => "00", 274 => "00", 275 => "00", 276 => "00", 277 => "00", 278 => "00", 279 => "00", 280 => "00", 281 => "00", 282 => "00", 283 => "00", 284 => "00", 285 => "00", 286 => "00", 287 => "00", 288 => "00", 289 => "00", 290 => "00", 291 => "00", 292 => "00", 293 => "00", 294 => "00", 295 => "00", 296 => "00", 297 => "00", 298 => "00", 299 => "00", 300 => "00", 301 => "00", 302 => "00", 303 => "00", 304 => "00", 305 => "00", 306 => "00", 307 => "00", 308 => "00", 309 => "00", 310 => "00", 311 => "00", 312 => "00", 313 => "00", 314 => "00", 315 => "00", 316 => "00", 317 => "00", 318 => "00", 319 => "00", 320 => "00", 321 => "00", 322 => "00", 323 => "00", 324 => "00", 325 => "00", 326 => "00", 327 => "00", 328 => "00", 329 => "00", 330 => "00", 331 => "00", 332 => "00", 333 => "00", 334 => "00", 335 => "00", 336 => "00", 337 => "00", 338 => "00", 339 => "00", 340 => "00", 341 => "00", 342 => "00", 343 => "00", 344 => "00", 345 => "00", 346 => "00", 347 => "00", 348 => "00", 349 => "00", 350 => "00", 351 => "00", 352 => "00", 353 => "00", 354 => "00", 355 => "00", 356 => "00", 357 => "00", 358 => "00", 359 => "00", 360 => "00", 361 => "00", 362 => "00", 363 => "00", 364 => "00", 365 => "00", 366 => "00", 367 => "00", 368 => "00", 369 => "00", 370 => "00", 371 => "00", 372 => "00", 373 => "00", 374 => "00", 375 => "00", 376 => "00", 377 => "00", 378 => "00", 379 => "00", 380 => "00", 381 => "00", 382 => "00", 383 => "00", 384 => "00", 385 => "00", 386 => "00", 387 => "00", 388 => "00", 389 => "00", 390 => "00", 391 => "00", 392 => "00", 393 => "00", 394 => "00", 395 => "00", 396 => "00", 397 => "00", 398 => "00", 399 => "00", 400 => "00", 401 => "00", 402 => "00", 403 => "00", 404 => "00", 405 => "00", 406 => "00", 407 => "00", 408 => "00", 409 => "00", 410 => "00", 411 => "00", 412 => "00", 413 => "00", 414 => "00", 415 => "00", 416 => "00", 417 => "00", 418 => "00", 419 => "00", 420 => "00", 421 => "00", 422 => "00", 423 => "00", 424 => "00", 425 => "00", 426 => "00", 427 => "00", 428 => "00", 429 => "00", 430 => "00", 431 => "00", 432 => "00", 433 => "00", 434 => "00", 435 => "00", 436 => "00", 437 => "00", 438 => "00", 439 => "00", 440 => "00", 441 => "00", 442 => "00", 443 => "00", 444 => "00", 445 => "00", 446 => "00", 447 => "00", 448 => "00", 449 => "00", 450 => "00", 451 => "00", 452 => "00", 453 => "00", 454 => "00", 455 => "00", 456 => "00", 457 => "00", 458 => "00", 459 => "00", 460 => "00", 461 => "00", 462 => "00", 463 => "00", 464 => "00", 465 => "00", 466 => "00", 467 => "00", 468 => "00", 469 => "00", 470 => "00", 471 => "00", 472 => "00", 473 => "00", 474 => "00", 475 => "00", 476 => "00", 477 => "00", 478 => "00", 479 => "00", 480 => "00", 481 => "00", 482 => "00", 483 => "00", 484 => "00", 485 => "00", 486 => "00", 487 => "00", 488 => "00", 489 => "00", 490 => "00", 491 => "00", 492 => "00", 493 => "00", 494 => "00", 495 => "00", 496 => "00", 497 => "00", 498 => "00", 499 => "00", 500 => "00", 501 => "00", 502 => "00", 503 => "00", 504 => "00", 505 => "00", 506 => "00", 507 => "00", 508 => "00", 509 => "00", 510 => "00", 511 => "00", 512 => "00", 513 => "00", 514 => "00", 515 => "00", 516 => "00", 517 => "00", 518 => "00", 519 => "00", 520 => "00", 521 => "00", 522 => "00", 523 => "00", 524 => "00", 525 => "00", 526 => "00", 527 => "00", 528 => "00", 529 => "00", 530 => "00", 531 => "00", 532 => "00", 533 => "00", 534 => "00", 535 => "00", 536 => "00", 537 => "00", 538 => "00", 539 => "00", 540 => "00", 541 => "00", 542 => "00", 543 => "00", 544 => "00", 545 => "00", 546 => "00", 547 => "00", 548 => "00", 549 => "00", 550 => "00", 551 => "00", 552 => "00", 553 => "00", 554 => "00", 555 => "00", 556 => "00", 557 => "00", 558 => "00", 559 => "00", 560 => "00", 561 => "00", 562 => "00", 563 => "00", 564 => "00", 565 => "00", 566 => "00", 567 => "00", 568 => "00", 569 => "00", 570 => "00", 571 => "00", 572 => "00", 573 => "00", 574 => "00", 575 => "00", 576 => "00", 577 => "00", 578 => "00", 579 => "00", 580 => "00", 581 => "00", 582 => "00", 583 => "00", 584 => "00", 585 => "00", 586 => "00", 587 => "00", 588 => "00", 589 => "00", 590 => "00", 591 => "00", 592 => "00", 593 => "00", 594 => "00", 595 => "00", 596 => "00", 597 => "00", 598 => "00", 599 => "00", 600 => "00", 601 => "00", 602 => "00", 603 => "00", 604 => "00", 605 => "00", 606 => "00", 607 => "00", 608 => "00", 609 => "00", 610 => "00", 611 => "00", 612 => "00", 613 => "00", 614 => "00", 615 => "00", 616 => "00", 617 => "00", 618 => "00", 619 => "00", 620 => "00", 621 => "00", 622 => "00", 623 => "00", 624 => "00", 625 => "00", 626 => "00", 627 => "00", 628 => "00", 629 => "00", 630 => "00", 631 => "00", 632 => "00", 633 => "00", 634 => "00", 635 => "00", 636 => "00", 637 => "00", 638 => "00", 639 => "00", 640 => "00", 641 => "00", 642 => "00", 643 => "00", 644 => "00", 645 => "00", 646 => "00", 647 => "00", 648 => "00", 649 => "00", 650 => "00", 651 => "00", 652 => "00", 653 => "00", 654 => "00", 655 => "00", 656 => "00", 657 => "00", 658 => "00", 659 => "00", 660 => "00", 661 => "00", 662 => "00", 663 => "00", 664 => "00", 665 => "00", 666 => "00", 667 => "00", 668 => "00", 669 => "00", 670 => "00", 671 => "00", 672 => "00", 673 => "00", 674 => "00", 675 => "00", 676 => "00", 677 => "00", 678 => "00", 679 => "00", 680 => "00", 681 => "00", 682 => "00", 683 => "00", 684 => "00", 685 => "00", 686 => "00", 687 => "00", 688 => "00", 689 => "00", 690 => "00", 691 => "00", 692 => "00", 693 => "00", 694 => "00", 695 => "00", 696 => "00", 697 => "00", 698 => "00", 699 => "00", 700 => "00", 701 => "00", 702 => "00", 703 => "00", 704 => "00", 705 => "00", 706 => "00", 707 => "00", 708 => "00", 709 => "00", 710 => "00", 711 => "00", 712 => "00", 713 => "00", 714 => "00", 715 => "00", 716 => "00", 717 => "00", 718 => "00", 719 => "00", 720 => "00", 721 => "00", 722 => "00", 723 => "00", 724 => "00", 725 => "00", 726 => "00", 727 => "00", 728 => "00", 729 => "00", 730 => "00", 731 => "00", 732 => "00", 733 => "00", 734 => "00", 735 => "00", 736 => "00", 737 => "00", 738 => "00", 739 => "00", 740 => "00", 741 => "00", 742 => "00", 743 => "00", 744 => "00", 745 => "00", 746 => "00", 747 => "00", 748 => "00", 749 => "00", 750 => "00", 751 => "00", 752 => "00", 753 => "00", 754 => "00", 755 => "00", 756 => "00", 757 => "00", 758 => "00", 759 => "00", 760 => "00", 761 => "00", 762 => "00", 763 => "00", 764 => "00", 765 => "00", 766 => "00", 767 => "00", 768 => "00", 769 => "00", 770 => "00", 771 => "00", 772 => "00", 773 => "00", 774 => "00", 775 => "00", 776 => "00", 777 => "00", 778 => "00", 779 => "00", 780 => "00", 781 => "00", 782 => "00", 783 => "00", 784 => "00", 785 => "00", 786 => "00", 787 => "00", 788 => "00", 789 => "00", 790 => "00", 791 => "00", 792 => "00", 793 => "00", 794 => "00", 795 => "00", 796 => "00", 797 => "00", 798 => "00", 799 => "00", 800 => "00", 801 => "00", 802 => "00", 803 => "00", 804 => "00", 805 => "00", 806 => "00", 807 => "00", 808 => "00", 809 => "00", 810 => "00", 811 => "00", 812 => "00", 813 => "00", 814 => "00", 815 => "00", 816 => "00", 817 => "00", 818 => "00", 819 => "00", 820 => "00", 821 => "00", 822 => "00", 823 => "00", 824 => "00", 825 => "00", 826 => "00", 827 => "00", 828 => "00", 829 => "00", 830 => "00", 831 => "00", 832 => "00", 833 => "00", 834 => "00", 835 => "00", 836 => "00", 837 => "00", 838 => "00", 839 => "00", 840 => "00", 841 => "00", 842 => "00", 843 => "00", 844 => "00", 845 => "00", 846 => "00", 847 => "00", 848 => "00", 849 => "00", 850 => "00", 851 => "00", 852 => "00", 853 => "00", 854 => "00", 855 => "00", 856 => "00", 857 => "00", 858 => "00", 859 => "00", 860 => "00", 861 => "00", 862 => "00", 863 => "00", 864 => "00", 865 => "00", 866 => "00", 867 => "00", 868 => "00", 869 => "00", 870 => "00", 871 => "00", 872 => "00", 873 => "00", 874 => "00", 875 => "00", 876 => "00", 877 => "00", 878 => "00", 879 => "00", 880 => "00", 881 => "00", 882 => "00", 883 => "00", 884 => "00", 885 => "00", 886 => "00", 887 => "00", 888 => "00", 889 => "00", 890 => "00", 891 => "00", 892 => "00", 893 => "00", 894 => "00", 895 => "00", 896 => "00", 897 => "00", 898 => "00", 899 => "00", 900 => "00", 901 => "00", 902 => "00", 903 => "00", 904 => "00", 905 => "00", 906 => "00", 907 => "00", 908 => "00", 909 => "00", 910 => "00", 911 => "00", 912 => "00", 913 => "00", 914 => "00", 915 => "00", 916 => "00", 917 => "00", 918 => "00", 919 => "00", 920 => "00", 921 => "00", 922 => "00", 923 => "00", 924 => "00", 925 => "00", 926 => "00", 927 => "00", 928 => "00", 929 => "00", 930 => "00", 931 => "00", 932 => "00", 933 => "00", 934 => "00", 935 => "00", 936 => "00", 937 => "00", 938 => "00", 939 => "00", 940 => "00", 941 => "00", 942 => "00", 943 => "00", 944 => "00", 945 => "00", 946 => "00", 947 => "00", 948 => "00", 949 => "00", 950 => "00", 951 => "00", 952 => "00", 953 => "00", 954 => "00", 955 => "00", 956 => "00", 957 => "00", 958 => "00", 959 => "00", 960 => "01", 961 => "11", 962 => "10", 963 => "11", 964 => "01", 965 => "11", 966 => "01", 967 => "00", 968 => "10", 969 => "11", 970 => "10", 971 => "11", 972 => "01", 973 => "11", 974 => "01", 975 => "00", 976 => "10", 977 => "11", 978 => "10", 979 => "11", 980 => "01", 981 => "11", 982 => "01", 983 => "00", 984 => "10", 985 => "11", 986 => "01", 987 => "00", 988 => "10", 989 => "00", 990 => "01", 991 => "11", 992 => "01", 993 => "00", 994 => "10", 995 => "00", 996 => "01", 997 => "00", 998 => "10", 999 => "00", 1000 => "01", 1001 => "11", 1002 => "10", 1003 => "00", 1004 => "01", 1005 => "11", 1006 => "01", 1007 => "11", 1008 => "10", 1009 => "00", 1010 => "01", 1011 => "11", 1012 => "10", 1013 => "00", 1014 => "10", 1015 => "11", 1016 => "01", 1017 => "00", 1018 => "10", 1019 => "00", 1020 => "01", 1021 => "11", 1022 => "10", 1023 => "00", 1024 => "10", 1025 => "11", 1026 => "01", 1027 => "00", 1028 => "10", 1029 => "00", 1030 => "01", 1031 => "11", 1032 => "10", 1033 => "00", 1034 => "10", 1035 => "11", 1036 => "10", 1037 => "11", 1038 => "01", 1039 => "11", 1040 => "10", 1041 => "00", 1042 => "10", 1043 => "11", 1044 => "10", 1045 => "11", 1046 => "01", 1047 => "11", 1048 => "01", 1049 => "00", 1050 => "10", 1051 => "11", 1052 => "10", 1053 => "11", 1054 => "01", 1055 => "11", 1056 => "01", 1057 => "00", 1058 => "10", 1059 => "11", 1060 => "10", 1061 => "11", 1062 => "01", 1063 => "11", 1064 => "01", 1065 => "00", 1066 => "00", 1067 => "00", 1068 => "00", 1069 => "00", 1070 => "00", 1071 => "00", 1072 => "00", 1073 => "00", 1074 => "00", 1075 => "00", 1076 => "00", 1077 => "00", 1078 => "00", 1079 => "00", 1080 => "00", 1081 => "00", 1082 => "00", 1083 => "00", 1084 => "00", 1085 => "00", 1086 => "00", 1087 => "00", 1088 => "00", 1089 => "00", 1090 => "00", 1091 => "00", 1092 => "00", 1093 => "00", 1094 => "00", 1095 => "00", 1096 => "00", 1097 => "00", 1098 => "00", 1099 => "00", 1100 => "00", 1101 => "00", 1102 => "00", 1103 => "00", 1104 => "00", 1105 => "00", 1106 => "00", 1107 => "00", 1108 => "00", 1109 => "00", 1110 => "00", 1111 => "00", 1112 => "00", 1113 => "00", 1114 => "00", 1115 => "00", 1116 => "00", 1117 => "00", 1118 => "00", 1119 => "00", 1120 => "00", 1121 => "00", 1122 => "00", 1123 => "00", 1124 => "00", 1125 => "00", 1126 => "00", 1127 => "00", 1128 => "00", 1129 => "00", 1130 => "00", 1131 => "00", 1132 => "00", 1133 => "00", 1134 => "00", 1135 => "00", 1136 => "00", 1137 => "00", 1138 => "00", 1139 => "00", 1140 => "00", 1141 => "00", 1142 => "00", 1143 => "00", 1144 => "00", 1145 => "00", 1146 => "00", 1147 => "00", 1148 => "00", 1149 => "00", 1150 => "00", 1151 => "00", 1152 => "00", 1153 => "00", 1154 => "00", 1155 => "00", 1156 => "00", 1157 => "00", 1158 => "00", 1159 => "00", 1160 => "00", 1161 => "00", 1162 => "00", 1163 => "00", 1164 => "00", 1165 => "00", 1166 => "00", 1167 => "00", 1168 => "00", 1169 => "00", 1170 => "00", 1171 => "00", 1172 => "00", 1173 => "00", 1174 => "00", 1175 => "00", 1176 => "00", 1177 => "00", 1178 => "00", 1179 => "00", 1180 => "00", 1181 => "00", 1182 => "00", 1183 => "00", 1184 => "00", 1185 => "00", 1186 => "00", 1187 => "00", 1188 => "00", 1189 => "00", 1190 => "00", 1191 => "00", 1192 => "00", 1193 => "00", 1194 => "00", 1195 => "00", 1196 => "00", 1197 => "00", 1198 => "00", 1199 => "00", 1200 => "00", 1201 => "00", 1202 => "00", 1203 => "00", 1204 => "00", 1205 => "00", 1206 => "00", 1207 => "00", 1208 => "00", 1209 => "00", 1210 => "00", 1211 => "00", 1212 => "00", 1213 => "00", 1214 => "00", 1215 => "00", 1216 => "00", 1217 => "00", 1218 => "00", 1219 => "00", 1220 => "00", 1221 => "00", 1222 => "00", 1223 => "00", 1224 => "00", 1225 => "00", 1226 => "00", 1227 => "00", 1228 => "00", 1229 => "00", 1230 => "00", 1231 => "00", 1232 => "00", 1233 => "00", 1234 => "00", 1235 => "00", 1236 => "00", 1237 => "00", 1238 => "00", 1239 => "00", 1240 => "00", 1241 => "00", 1242 => "00", 1243 => "00", 1244 => "00", 1245 => "00", 1246 => "00", 1247 => "00", 1248 => "00", 1249 => "00", 1250 => "00", 1251 => "00", 1252 => "00", 1253 => "00", 1254 => "00", 1255 => "00", 1256 => "00", 1257 => "00", 1258 => "00", 1259 => "00", 1260 => "00", 1261 => "00", 1262 => "00", 1263 => "00", 1264 => "00", 1265 => "00", 1266 => "00", 1267 => "00", 1268 => "00", 1269 => "00", 1270 => "00", 1271 => "00", 1272 => "00", 1273 => "00", 1274 => "00", 1275 => "00", 1276 => "00", 1277 => "00", 1278 => "00", 1279 => "00", 1280 => "00", 1281 => "00", 1282 => "00", 1283 => "00", 1284 => "00", 1285 => "00", 1286 => "00", 1287 => "00", 1288 => "00", 1289 => "00", 1290 => "00", 1291 => "00", 1292 => "00", 1293 => "00", 1294 => "00", 1295 => "00", 1296 => "00", 1297 => "00", 1298 => "00", 1299 => "00", 1300 => "00", 1301 => "00", 1302 => "00", 1303 => "00", 1304 => "00", 1305 => "00", 1306 => "00", 1307 => "00", 1308 => "00", 1309 => "00", 1310 => "00", 1311 => "00", 1312 => "00", 1313 => "00", 1314 => "00", 1315 => "00", 1316 => "00", 1317 => "00", 1318 => "00", 1319 => "00", 1320 => "00", 1321 => "00", 1322 => "00", 1323 => "00", 1324 => "00", 1325 => "00", 1326 => "00", 1327 => "00", 1328 => "00", 1329 => "00", 1330 => "00", 1331 => "00", 1332 => "00", 1333 => "00", 1334 => "00", 1335 => "00", 1336 => "00", 1337 => "00", 1338 => "00", 1339 => "00", 1340 => "00", 1341 => "00", 1342 => "00", 1343 => "00", 1344 => "00", 1345 => "00", 1346 => "00", 1347 => "00", 1348 => "00", 1349 => "00", 1350 => "00", 1351 => "00", 1352 => "00", 1353 => "00", 1354 => "00", 1355 => "00", 1356 => "00", 1357 => "00", 1358 => "00", 1359 => "00", 1360 => "00", 1361 => "00", 1362 => "00", 1363 => "00", 1364 => "00", 1365 => "00", 1366 => "00", 1367 => "00", 1368 => "00", 1369 => "00", 1370 => "00", 1371 => "00", 1372 => "00", 1373 => "00", 1374 => "00", 1375 => "00", 1376 => "00", 1377 => "00", 1378 => "00", 1379 => "00", 1380 => "00", 1381 => "00", 1382 => "00", 1383 => "00", 1384 => "00", 1385 => "00", 1386 => "00", 1387 => "00", 1388 => "00", 1389 => "00", 1390 => "00", 1391 => "00", 1392 => "00", 1393 => "00", 1394 => "00", 1395 => "00", 1396 => "00", 1397 => "00", 1398 => "00", 1399 => "00", 1400 => "00", 1401 => "00", 1402 => "00", 1403 => "00", 1404 => "00", 1405 => "00", 1406 => "00", 1407 => "00", 1408 => "00", 1409 => "00", 1410 => "00", 1411 => "00", 1412 => "00", 1413 => "00", 1414 => "00", 1415 => "00", 1416 => "00", 1417 => "00", 1418 => "00", 1419 => "00", 1420 => "00", 1421 => "00", 1422 => "00", 1423 => "00", 1424 => "00", 1425 => "00", 1426 => "00", 1427 => "00", 1428 => "00", 1429 => "00", 1430 => "00", 1431 => "00", 1432 => "00", 1433 => "00", 1434 => "00", 1435 => "00", 1436 => "00", 1437 => "00", 1438 => "00", 1439 => "00", 1440 => "00", 1441 => "00", 1442 => "00", 1443 => "00", 1444 => "00", 1445 => "00", 1446 => "00", 1447 => "00", 1448 => "00", 1449 => "00", 1450 => "00", 1451 => "00", 1452 => "00", 1453 => "00", 1454 => "00", 1455 => "00", 1456 => "00", 1457 => "00", 1458 => "00", 1459 => "00", 1460 => "00", 1461 => "00", 1462 => "00", 1463 => "00", 1464 => "00", 1465 => "00", 1466 => "00", 1467 => "00", 1468 => "00", 1469 => "00", 1470 => "00", 1471 => "00", 1472 => "00", 1473 => "00", 1474 => "00", 1475 => "00", 1476 => "00", 1477 => "00", 1478 => "00", 1479 => "00", 1480 => "00", 1481 => "00", 1482 => "00", 1483 => "00", 1484 => "00", 1485 => "00", 1486 => "00", 1487 => "00", 1488 => "00", 1489 => "00", 1490 => "00", 1491 => "00", 1492 => "00", 1493 => "00", 1494 => "00", 1495 => "00", 1496 => "00", 1497 => "00", 1498 => "00", 1499 => "00", 1500 => "00", 1501 => "00", 1502 => "00", 1503 => "00", 1504 => "00", 1505 => "00", 1506 => "00", 1507 => "00", 1508 => "00", 1509 => "00", 1510 => "00", 1511 => "00", 1512 => "00", 1513 => "00", 1514 => "00", 1515 => "00", 1516 => "00", 1517 => "00", 1518 => "00", 1519 => "00", 1520 => "00", 1521 => "00", 1522 => "00", 1523 => "00", 1524 => "00", 1525 => "00", 1526 => "00", 1527 => "00", 1528 => "00", 1529 => "00", 1530 => "00", 1531 => "00", 1532 => "00", 1533 => "00", 1534 => "00", 1535 => "00", 1536 => "00", 1537 => "00", 1538 => "00", 1539 => "00", 1540 => "00", 1541 => "00", 1542 => "00", 1543 => "00", 1544 => "00", 1545 => "00", 1546 => "00", 1547 => "00", 1548 => "00", 1549 => "00", 1550 => "00", 1551 => "00", 1552 => "00", 1553 => "00", 1554 => "00", 1555 => "00", 1556 => "00", 1557 => "00", 1558 => "00", 1559 => "00", 1560 => "00", 1561 => "00", 1562 => "00", 1563 => "00", 1564 => "00", 1565 => "00", 1566 => "00", 1567 => "00", 1568 => "00", 1569 => "00", 1570 => "00", 1571 => "00", 1572 => "00", 1573 => "00", 1574 => "00", 1575 => "00", 1576 => "00", 1577 => "00", 1578 => "00", 1579 => "00", 1580 => "00", 1581 => "00", 1582 => "00", 1583 => "00", 1584 => "00", 1585 => "00", 1586 => "00", 1587 => "00", 1588 => "00", 1589 => "00", 1590 => "00", 1591 => "00", 1592 => "00", 1593 => "00", 1594 => "00", 1595 => "00", 1596 => "00", 1597 => "00", 1598 => "00", 1599 => "00", 1600 => "00", 1601 => "00", 1602 => "00", 1603 => "00", 1604 => "00", 1605 => "00", 1606 => "00", 1607 => "00", 1608 => "00", 1609 => "00", 1610 => "00", 1611 => "00", 1612 => "00", 1613 => "00", 1614 => "00", 1615 => "00", 1616 => "00", 1617 => "00", 1618 => "00", 1619 => "00", 1620 => "00", 1621 => "00", 1622 => "00", 1623 => "00", 1624 => "00", 1625 => "00", 1626 => "00", 1627 => "00", 1628 => "00", 1629 => "00", 1630 => "00", 1631 => "00", 1632 => "00", 1633 => "00", 1634 => "00", 1635 => "00", 1636 => "00", 1637 => "00", 1638 => "00", 1639 => "00", 1640 => "00", 1641 => "00", 1642 => "00", 1643 => "00", 1644 => "00", 1645 => "00", 1646 => "00", 1647 => "00", 1648 => "00", 1649 => "00", 1650 => "00", 1651 => "00", 1652 => "00", 1653 => "00", 1654 => "00", 1655 => "00", 1656 => "00", 1657 => "00", 1658 => "00", 1659 => "00", 1660 => "00", 1661 => "00", 1662 => "00", 1663 => "00", 1664 => "00", 1665 => "00", 1666 => "00", 1667 => "00", 1668 => "00", 1669 => "00", 1670 => "00", 1671 => "00", 1672 => "00", 1673 => "00", 1674 => "00", 1675 => "00", 1676 => "00", 1677 => "00", 1678 => "00", 1679 => "00", 1680 => "00", 1681 => "00", 1682 => "00", 1683 => "00", 1684 => "00", 1685 => "00", 1686 => "00", 1687 => "00", 1688 => "00", 1689 => "00", 1690 => "00", 1691 => "00", 1692 => "00", 1693 => "00", 1694 => "00", 1695 => "00", 1696 => "00", 1697 => "00", 1698 => "00", 1699 => "00", 1700 => "00", 1701 => "00", 1702 => "00", 1703 => "00", 1704 => "00", 1705 => "00", 1706 => "00", 1707 => "00", 1708 => "00", 1709 => "00", 1710 => "00", 1711 => "00", 1712 => "00", 1713 => "00", 1714 => "00", 1715 => "00", 1716 => "00", 1717 => "00", 1718 => "00", 1719 => "00", 1720 => "00", 1721 => "00", 1722 => "00", 1723 => "00", 1724 => "00", 1725 => "00", 1726 => "00", 1727 => "00", 1728 => "00", 1729 => "00", 1730 => "00", 1731 => "00", 1732 => "00", 1733 => "00", 1734 => "00", 1735 => "00", 1736 => "00", 1737 => "00", 1738 => "00", 1739 => "00", 1740 => "00", 1741 => "00", 1742 => "00", 1743 => "00", 1744 => "00", 1745 => "00", 1746 => "00", 1747 => "00", 1748 => "00", 1749 => "00", 1750 => "00", 1751 => "00", 1752 => "00", 1753 => "00", 1754 => "00", 1755 => "00", 1756 => "00", 1757 => "00", 1758 => "00", 1759 => "00", 1760 => "00", 1761 => "00", 1762 => "00", 1763 => "00", 1764 => "00", 1765 => "00", 1766 => "00", 1767 => "00", 1768 => "00", 1769 => "00", 1770 => "00", 1771 => "00", 1772 => "00", 1773 => "00", 1774 => "00", 1775 => "00", 1776 => "00", 1777 => "00", 1778 => "00", 1779 => "00", 1780 => "00", 1781 => "00", 1782 => "00", 1783 => "00", 1784 => "00", 1785 => "00", 1786 => "00", 1787 => "00", 1788 => "00", 1789 => "00", 1790 => "00", 1791 => "00", 1792 => "00", 1793 => "00", 1794 => "00", 1795 => "00", 1796 => "00", 1797 => "00", 1798 => "00", 1799 => "00", 1800 => "00", 1801 => "00", 1802 => "00", 1803 => "00", 1804 => "00", 1805 => "00", 1806 => "00", 1807 => "00", 1808 => "00", 1809 => "00", 1810 => "00", 1811 => "00", 1812 => "00", 1813 => "00", 1814 => "00", 1815 => "00", 1816 => "00", 1817 => "00", 1818 => "00", 1819 => "00", 1820 => "00", 1821 => "00", 1822 => "00", 1823 => "00", 1824 => "00", 1825 => "00", 1826 => "00", 1827 => "00", 1828 => "00", 1829 => "00", 1830 => "00", 1831 => "00", 1832 => "00", 1833 => "00", 1834 => "00", 1835 => "00", 1836 => "00", 1837 => "00", 1838 => "00", 1839 => "00", 1840 => "00", 1841 => "00", 1842 => "00", 1843 => "00", 1844 => "00", 1845 => "00", 1846 => "00", 1847 => "00", 1848 => "00", 1849 => "00", 1850 => "00", 1851 => "00", 1852 => "00", 1853 => "00", 1854 => "00", 1855 => "00", 1856 => "00", 1857 => "00", 1858 => "00", 1859 => "00", 1860 => "00", 1861 => "00", 1862 => "00", 1863 => "00", 1864 => "00", 1865 => "00", 1866 => "00", 1867 => "00", 1868 => "00", 1869 => "00", 1870 => "00", 1871 => "00", 1872 => "00", 1873 => "00", 1874 => "00", 1875 => "00", 1876 => "00", 1877 => "00", 1878 => "00", 1879 => "00", 1880 => "00", 1881 => "00", 1882 => "00", 1883 => "00", 1884 => "00", 1885 => "00", 1886 => "00", 1887 => "00", 1888 => "00", 1889 => "00", 1890 => "00", 1891 => "00", 1892 => "00", 1893 => "00", 1894 => "00", 1895 => "00", 1896 => "00", 1897 => "00", 1898 => "00", 1899 => "00", 1900 => "00", 1901 => "00", 1902 => "00", 1903 => "00", 1904 => "00", 1905 => "00", 1906 => "00", 1907 => "00", 1908 => "00", 1909 => "00", 1910 => "00", 1911 => "00", 1912 => "00", 1913 => "00", 1914 => "00", 1915 => "00", 1916 => "00", 1917 => "00", 1918 => "00", 1919 => "00", 1920 => "00", 1921 => "00", 1922 => "00", 1923 => "00", 1924 => "00", 1925 => "00", 1926 => "00", 1927 => "00", 1928 => "00", 1929 => "00", 1930 => "00", 1931 => "00", 1932 => "00", 1933 => "00", 1934 => "00", 1935 => "00", 1936 => "00", 1937 => "00", 1938 => "00", 1939 => "00", 1940 => "00", 1941 => "00", 1942 => "00", 1943 => "00", 1944 => "00", 1945 => "00", 1946 => "00", 1947 => "00", 1948 => "00", 1949 => "00", 1950 => "00", 1951 => "00", 1952 => "00", 1953 => "00", 1954 => "00", 1955 => "00", 1956 => "00", 1957 => "00", 1958 => "00", 1959 => "00", 1960 => "00", 1961 => "00", 1962 => "00", 1963 => "00", 1964 => "00", 1965 => "00", 1966 => "00", 1967 => "00", 1968 => "00", 1969 => "00", 1970 => "00", 1971 => "00", 1972 => "00", 1973 => "00", 1974 => "00", 1975 => "00", 1976 => "00", 1977 => "00", 1978 => "00", 1979 => "00", 1980 => "00", 1981 => "00", 1982 => "00", 1983 => "00", 1984 => "00", 1985 => "00", 1986 => "00", 1987 => "00", 1988 => "00", 1989 => "00", 1990 => "00", 1991 => "00", 1992 => "00", 1993 => "00", 1994 => "00", 1995 => "00", 1996 => "00", 1997 => "00", 1998 => "00", 1999 => "00", 2000 => "00", 2001 => "00", 2002 => "00", 2003 => "00", 2004 => "00", 2005 => "00", 2006 => "00", 2007 => "00", 2008 => "00", 2009 => "00", 2010 => "00", 2011 => "00", 2012 => "00", 2013 => "00", 2014 => "00", 2015 => "00", 2016 => "00", 2017 => "00", 2018 => "00", 2019 => "00", 2020 => "00", 2021 => "00", 2022 => "00", 2023 => "00", 2024 => "00", 2025 => "00", 2026 => "01", 2027 => "11", 2028 => "10", 2029 => "11", 2030 => "01", 2031 => "11", 2032 => "01", 2033 => "00", 2034 => "10", 2035 => "11", 2036 => "10", 2037 => "11", 2038 => "01", 2039 => "11", 2040 => "01", 2041 => "00", 2042 => "10", 2043 => "11", 2044 => "10", 2045 => "11", 2046 => "01", 2047 => "11", 2048 => "01", 2049 => "00", 2050 => "10", 2051 => "11", 2052 => "10", 2053 => "11", 2054 => "01", 2055 => "11", 2056 => "01", 2057 => "00", 2058 => "10", 2059 => "11", 2060 => "10", 2061 => "11", 2062 => "01", 2063 => "11", 2064 => "01", 2065 => "00", 2066 => "10", 2067 => "11", 2068 => "10", 2069 => "11", 2070 => "01", 2071 => "11", 2072 => "01", 2073 => "00", 2074 => "10", 2075 => "11", 2076 => "10", 2077 => "11", 2078 => "01", 2079 => "11", 2080 => "01", 2081 => "00", 2082 => "10", 2083 => "11", 2084 => "10", 2085 => "11", 2086 => "01", 2087 => "11", 2088 => "01", 2089 => "00", 2090 => "10", 2091 => "11", 2092 => "10", 2093 => "11", 2094 => "01", 2095 => "11", 2096 => "01", 2097 => "00", 2098 => "10", 2099 => "11", 2100 => "10", 2101 => "11", 2102 => "01", 2103 => "11", 2104 => "01", 2105 => "00", 2106 => "10", 2107 => "11", 2108 => "10", 2109 => "11", 2110 => "01", 2111 => "11", 2112 => "01", 2113 => "00", 2114 => "10", 2115 => "11", 2116 => "10", 2117 => "11", 2118 => "01", 2119 => "11", 2120 => "01", 2121 => "00", 2122 => "10", 2123 => "11", 2124 => "10", 2125 => "11", 2126 => "01", 2127 => "11", 2128 => "01", 2129 => "00", 2130 => "10", 2131 => "11", 2132 => "10", 2133 => "11", 2134 => "01", 2135 => "11", 2136 => "01", 2137 => "00", 2138 => "10", 2139 => "11", 2140 => "10", 2141 => "11", 2142 => "01", 2143 => "11", 2144 => "01", 2145 => "00", 2146 => "10", 2147 => "11", 2148 => "10", 2149 => "11", 2150 => "01", 2151 => "11", 2152 => "01", 2153 => "00", 2154 => "10", 2155 => "11", 2156 => "10", 2157 => "11", 2158 => "01", 2159 => "11", 2160 => "01", 2161 => "00", 2162 => "10", 2163 => "11", 2164 => "10", 2165 => "11", 2166 => "01", 2167 => "11", 2168 => "01", 2169 => "00", 2170 => "10", 2171 => "11", 2172 => "01", 2173 => "00", 2174 => "00", 2175 => "00", 2176 => "00", 2177 => "00", 2178 => "00", 2179 => "00", 2180 => "00", 2181 => "00", 2182 => "00", 2183 => "00", 2184 => "00", 2185 => "00", 2186 => "00", 2187 => "00", 2188 => "00", 2189 => "00", 2190 => "00", 2191 => "00", 2192 => "00", 2193 => "00", 2194 => "00", 2195 => "00", 2196 => "00", 2197 => "00", 2198 => "00", 2199 => "00", 2200 => "00", 2201 => "00", 2202 => "00", 2203 => "00", 2204 => "00", 2205 => "00", 2206 => "00", 2207 => "00", 2208 => "00", 2209 => "00", 2210 => "00", 2211 => "00", 2212 => "00", 2213 => "00", 2214 => "00", 2215 => "00", 2216 => "00", 2217 => "00", 2218 => "00", 2219 => "00", 2220 => "00", 2221 => "00", 2222 => "00", 2223 => "00", 2224 => "00", 2225 => "00", 2226 => "00", 2227 => "00", 2228 => "00", 2229 => "00", 2230 => "00", 2231 => "00", 2232 => "00", 2233 => "00", 2234 => "00", 2235 => "00", 2236 => "00", 2237 => "00", 2238 => "00", 2239 => "00", 2240 => "00", 2241 => "00", 2242 => "00", 2243 => "00", 2244 => "00", 2245 => "00", 2246 => "00", 2247 => "00", 2248 => "00", 2249 => "00", 2250 => "00", 2251 => "00", 2252 => "00", 2253 => "00", 2254 => "00", 2255 => "00", 2256 => "00", 2257 => "00", 2258 => "00", 2259 => "00", 2260 => "00", 2261 => "00", 2262 => "00", 2263 => "00", 2264 => "00", 2265 => "00", 2266 => "00", 2267 => "00", 2268 => "00", 2269 => "00", 2270 => "00", 2271 => "00", 2272 => "00", 2273 => "00", 2274 => "00", 2275 => "00", 2276 => "00", 2277 => "00", 2278 => "00", 2279 => "00", 2280 => "00", 2281 => "00", 2282 => "00", 2283 => "00", 2284 => "00", 2285 => "00", 2286 => "00", 2287 => "00", 2288 => "00", 2289 => "00", 2290 => "00", 2291 => "00", 2292 => "00", 2293 => "00", 2294 => "00", 2295 => "00", 2296 => "00", 2297 => "00", 2298 => "00", 2299 => "00", 2300 => "00", 2301 => "00", 2302 => "00", 2303 => "00", 2304 => "00", 2305 => "00", 2306 => "00", 2307 => "00", 2308 => "00", 2309 => "00", 2310 => "00", 2311 => "00", 2312 => "00", 2313 => "00", 2314 => "00", 2315 => "00", 2316 => "00", 2317 => "00", 2318 => "00", 2319 => "00", 2320 => "00", 2321 => "00", 2322 => "00", 2323 => "00", 2324 => "00", 2325 => "00", 2326 => "00", 2327 => "00", 2328 => "00", 2329 => "00", 2330 => "00", 2331 => "00", 2332 => "00", 2333 => "00", 2334 => "00", 2335 => "00", 2336 => "00", 2337 => "00", 2338 => "00", 2339 => "00", 2340 => "00", 2341 => "00", 2342 => "00", 2343 => "00", 2344 => "00", 2345 => "00", 2346 => "00", 2347 => "00", 2348 => "00", 2349 => "00", 2350 => "00", 2351 => "00", 2352 => "00", 2353 => "00", 2354 => "00", 2355 => "00", 2356 => "00", 2357 => "00", 2358 => "00", 2359 => "00", 2360 => "00", 2361 => "00", 2362 => "00", 2363 => "00", 2364 => "00", 2365 => "00", 2366 => "00", 2367 => "00", 2368 => "00", 2369 => "00", 2370 => "00", 2371 => "00", 2372 => "00", 2373 => "00", 2374 => "00", 2375 => "00", 2376 => "00", 2377 => "00", 2378 => "00", 2379 => "00", 2380 => "00", 2381 => "00", 2382 => "00", 2383 => "00", 2384 => "00", 2385 => "00", 2386 => "00", 2387 => "00", 2388 => "00", 2389 => "00", 2390 => "00", 2391 => "00", 2392 => "00", 2393 => "00", 2394 => "00", 2395 => "00", 2396 => "00", 2397 => "00", 2398 => "00", 2399 => "00", 2400 => "00", 2401 => "00", 2402 => "00", 2403 => "00", 2404 => "00", 2405 => "00", 2406 => "00", 2407 => "00", 2408 => "00", 2409 => "00", 2410 => "00", 2411 => "00", 2412 => "00", 2413 => "00", 2414 => "00", 2415 => "00", 2416 => "00", 2417 => "00", 2418 => "00", 2419 => "00", 2420 => "00", 2421 => "00", 2422 => "00", 2423 => "00", 2424 => "00", 2425 => "00", 2426 => "00", 2427 => "00", 2428 => "00", 2429 => "00", 2430 => "00", 2431 => "00", 2432 => "00", 2433 => "00", 2434 => "00", 2435 => "00", 2436 => "00", 2437 => "00", 2438 => "00", 2439 => "00", 2440 => "00", 2441 => "00", 2442 => "00", 2443 => "00", 2444 => "00", 2445 => "00", 2446 => "00", 2447 => "00", 2448 => "00", 2449 => "00", 2450 => "00", 2451 => "00", 2452 => "00", 2453 => "00", 2454 => "00", 2455 => "00", 2456 => "00", 2457 => "00", 2458 => "00", 2459 => "00", 2460 => "00", 2461 => "00", 2462 => "00", 2463 => "00", 2464 => "00", 2465 => "00", 2466 => "00", 2467 => "00", 2468 => "00", 2469 => "00", 2470 => "00", 2471 => "00", 2472 => "00", 2473 => "00", 2474 => "00", 2475 => "00", 2476 => "00", 2477 => "00", 2478 => "00", 2479 => "00", 2480 => "00", 2481 => "00", 2482 => "00", 2483 => "00", 2484 => "00", 2485 => "00", 2486 => "00", 2487 => "00", 2488 => "00", 2489 => "00", 2490 => "00", 2491 => "00", 2492 => "00", 2493 => "00", 2494 => "00", 2495 => "00", 2496 => "00", 2497 => "00", 2498 => "00", 2499 => "00", 2500 => "00", 2501 => "00", 2502 => "00", 2503 => "00", 2504 => "00", 2505 => "00", 2506 => "00", 2507 => "00", 2508 => "00", 2509 => "00", 2510 => "00", 2511 => "00", 2512 => "00", 2513 => "00", 2514 => "00", 2515 => "00", 2516 => "00", 2517 => "00", 2518 => "00", 2519 => "00", 2520 => "00", 2521 => "00", 2522 => "00", 2523 => "00", 2524 => "00", 2525 => "00", 2526 => "00", 2527 => "00", 2528 => "00", 2529 => "00", 2530 => "00", 2531 => "00", 2532 => "00", 2533 => "00", 2534 => "00", 2535 => "00", 2536 => "00", 2537 => "00", 2538 => "00", 2539 => "00", 2540 => "00", 2541 => "00", 2542 => "00", 2543 => "00", 2544 => "00", 2545 => "00", 2546 => "00", 2547 => "00", 2548 => "00", 2549 => "00", 2550 => "00", 2551 => "00", 2552 => "00", 2553 => "00", 2554 => "00", 2555 => "00", 2556 => "00", 2557 => "00", 2558 => "00", 2559 => "00", 2560 => "00", 2561 => "00", 2562 => "00", 2563 => "00", 2564 => "00", 2565 => "00", 2566 => "00", 2567 => "00", 2568 => "00", 2569 => "00", 2570 => "00", 2571 => "00", 2572 => "00", 2573 => "00", 2574 => "00", 2575 => "00", 2576 => "00", 2577 => "00", 2578 => "00", 2579 => "00", 2580 => "00", 2581 => "00", 2582 => "00", 2583 => "00", 2584 => "00", 2585 => "00", 2586 => "00", 2587 => "00", 2588 => "00", 2589 => "00", 2590 => "00", 2591 => "00", 2592 => "00", 2593 => "00", 2594 => "00", 2595 => "00", 2596 => "00", 2597 => "00", 2598 => "00", 2599 => "00", 2600 => "00", 2601 => "00", 2602 => "00", 2603 => "00", 2604 => "00", 2605 => "00", 2606 => "00", 2607 => "00", 2608 => "00", 2609 => "00", 2610 => "00", 2611 => "00", 2612 => "00", 2613 => "00", 2614 => "00", 2615 => "00", 2616 => "00", 2617 => "00", 2618 => "00", 2619 => "00", 2620 => "00", 2621 => "00", 2622 => "00", 2623 => "00", 2624 => "00", 2625 => "00", 2626 => "00", 2627 => "00", 2628 => "00", 2629 => "00", 2630 => "00", 2631 => "00", 2632 => "00", 2633 => "00", 2634 => "00", 2635 => "00", 2636 => "00", 2637 => "00", 2638 => "00", 2639 => "00", 2640 => "00", 2641 => "00", 2642 => "00", 2643 => "00", 2644 => "00", 2645 => "00", 2646 => "00", 2647 => "00", 2648 => "00", 2649 => "00", 2650 => "00", 2651 => "00", 2652 => "00", 2653 => "00", 2654 => "00", 2655 => "00", 2656 => "00", 2657 => "00", 2658 => "00", 2659 => "00", 2660 => "00", 2661 => "00", 2662 => "00", 2663 => "00", 2664 => "00", 2665 => "00", 2666 => "00", 2667 => "00", 2668 => "00", 2669 => "00", 2670 => "00", 2671 => "00", 2672 => "00", 2673 => "00", 2674 => "00", 2675 => "00", 2676 => "00", 2677 => "00", 2678 => "00", 2679 => "00", 2680 => "00", 2681 => "00", 2682 => "00", 2683 => "00", 2684 => "00", 2685 => "00", 2686 => "00", 2687 => "00", 2688 => "00", 2689 => "00", 2690 => "00", 2691 => "00", 2692 => "00", 2693 => "00", 2694 => "00", 2695 => "00", 2696 => "00", 2697 => "00", 2698 => "00", 2699 => "00", 2700 => "00", 2701 => "00", 2702 => "00", 2703 => "00", 2704 => "00", 2705 => "00", 2706 => "00", 2707 => "00", 2708 => "00", 2709 => "00", 2710 => "00", 2711 => "00", 2712 => "00", 2713 => "00", 2714 => "00", 2715 => "00", 2716 => "00", 2717 => "00", 2718 => "00", 2719 => "00", 2720 => "00", 2721 => "00", 2722 => "00", 2723 => "00", 2724 => "00", 2725 => "00", 2726 => "00", 2727 => "00", 2728 => "00", 2729 => "00", 2730 => "00", 2731 => "00", 2732 => "00", 2733 => "00", 2734 => "00", 2735 => "00", 2736 => "00", 2737 => "00", 2738 => "00", 2739 => "00", 2740 => "00", 2741 => "00", 2742 => "00", 2743 => "00", 2744 => "00", 2745 => "00", 2746 => "00", 2747 => "00", 2748 => "00", 2749 => "00", 2750 => "00", 2751 => "00", 2752 => "00", 2753 => "00", 2754 => "00", 2755 => "00", 2756 => "00", 2757 => "00", 2758 => "00", 2759 => "00", 2760 => "00", 2761 => "00", 2762 => "00", 2763 => "00", 2764 => "00", 2765 => "00", 2766 => "00", 2767 => "00", 2768 => "00", 2769 => "00", 2770 => "00", 2771 => "00", 2772 => "00", 2773 => "00", 2774 => "00", 2775 => "00", 2776 => "00", 2777 => "00", 2778 => "00", 2779 => "00", 2780 => "00", 2781 => "00", 2782 => "00", 2783 => "00", 2784 => "00", 2785 => "00", 2786 => "00", 2787 => "00", 2788 => "00", 2789 => "00", 2790 => "00", 2791 => "00", 2792 => "00", 2793 => "00", 2794 => "00", 2795 => "00", 2796 => "00", 2797 => "00", 2798 => "00", 2799 => "00", 2800 => "00", 2801 => "00", 2802 => "00", 2803 => "00", 2804 => "00", 2805 => "00", 2806 => "00", 2807 => "00", 2808 => "00", 2809 => "00", 2810 => "00", 2811 => "00", 2812 => "00", 2813 => "00", 2814 => "00", 2815 => "00", 2816 => "00", 2817 => "00", 2818 => "00", 2819 => "00", 2820 => "00", 2821 => "00", 2822 => "00", 2823 => "00", 2824 => "00", 2825 => "00", 2826 => "00", 2827 => "00", 2828 => "00", 2829 => "00", 2830 => "00", 2831 => "00", 2832 => "00", 2833 => "00", 2834 => "00", 2835 => "00", 2836 => "00", 2837 => "00", 2838 => "00", 2839 => "00", 2840 => "00", 2841 => "00", 2842 => "00", 2843 => "00", 2844 => "00", 2845 => "00", 2846 => "00", 2847 => "00", 2848 => "00", 2849 => "00", 2850 => "00", 2851 => "00", 2852 => "00", 2853 => "00", 2854 => "00", 2855 => "00", 2856 => "00", 2857 => "00", 2858 => "00", 2859 => "00", 2860 => "00", 2861 => "00", 2862 => "00", 2863 => "00", 2864 => "00", 2865 => "00", 2866 => "00", 2867 => "00", 2868 => "00", 2869 => "00", 2870 => "00", 2871 => "00", 2872 => "00", 2873 => "00", 2874 => "00", 2875 => "00", 2876 => "00", 2877 => "00", 2878 => "00", 2879 => "00", 2880 => "00", 2881 => "00", 2882 => "00", 2883 => "00", 2884 => "00", 2885 => "00", 2886 => "00", 2887 => "00", 2888 => "00", 2889 => "00", 2890 => "00", 2891 => "00", 2892 => "00", 2893 => "00", 2894 => "00", 2895 => "00", 2896 => "00", 2897 => "00", 2898 => "00", 2899 => "00", 2900 => "00", 2901 => "00", 2902 => "00", 2903 => "00", 2904 => "00", 2905 => "00", 2906 => "00", 2907 => "00", 2908 => "00", 2909 => "00", 2910 => "00", 2911 => "00", 2912 => "00", 2913 => "00", 2914 => "00", 2915 => "00", 2916 => "00", 2917 => "00", 2918 => "00", 2919 => "00", 2920 => "00", 2921 => "00", 2922 => "00", 2923 => "00", 2924 => "00", 2925 => "00", 2926 => "00", 2927 => "00", 2928 => "00", 2929 => "00", 2930 => "00", 2931 => "00", 2932 => "00", 2933 => "00", 2934 => "00", 2935 => "00", 2936 => "00", 2937 => "00", 2938 => "00", 2939 => "00", 2940 => "00", 2941 => "00", 2942 => "00", 2943 => "00", 2944 => "00", 2945 => "00", 2946 => "00", 2947 => "00", 2948 => "00", 2949 => "00", 2950 => "00", 2951 => "00", 2952 => "00", 2953 => "00", 2954 => "00", 2955 => "00", 2956 => "00", 2957 => "00", 2958 => "00", 2959 => "00", 2960 => "00", 2961 => "00", 2962 => "00", 2963 => "00", 2964 => "00", 2965 => "00", 2966 => "00", 2967 => "00", 2968 => "00", 2969 => "00", 2970 => "00", 2971 => "00", 2972 => "00", 2973 => "00", 2974 => "00", 2975 => "00", 2976 => "00", 2977 => "00", 2978 => "00", 2979 => "00", 2980 => "00", 2981 => "00", 2982 => "00", 2983 => "00", 2984 => "00", 2985 => "00", 2986 => "00", 2987 => "00", 2988 => "00", 2989 => "00", 2990 => "00", 2991 => "00", 2992 => "00", 2993 => "00", 2994 => "00", 2995 => "00", 2996 => "00", 2997 => "00", 2998 => "00", 2999 => "00", 3000 => "00", 3001 => "00", 3002 => "00", 3003 => "00", 3004 => "00", 3005 => "00", 3006 => "00", 3007 => "00", 3008 => "00", 3009 => "00", 3010 => "00", 3011 => "00", 3012 => "00", 3013 => "00", 3014 => "00", 3015 => "00", 3016 => "00", 3017 => "00", 3018 => "00", 3019 => "00", 3020 => "00", 3021 => "00", 3022 => "00", 3023 => "00", 3024 => "00", 3025 => "00", 3026 => "00", 3027 => "00", 3028 => "00", 3029 => "00", 3030 => "00", 3031 => "00", 3032 => "00", 3033 => "00", 3034 => "00", 3035 => "00", 3036 => "00", 3037 => "00", 3038 => "00", 3039 => "00", 3040 => "00", 3041 => "00", 3042 => "00", 3043 => "00", 3044 => "00", 3045 => "00", 3046 => "00", 3047 => "00", 3048 => "00", 3049 => "00", 3050 => "00", 3051 => "00", 3052 => "00", 3053 => "00", 3054 => "00", 3055 => "00", 3056 => "00", 3057 => "00", 3058 => "00", 3059 => "00", 3060 => "00", 3061 => "00", 3062 => "00", 3063 => "00", 3064 => "00", 3065 => "00", 3066 => "00", 3067 => "00", 3068 => "00", 3069 => "00", 3070 => "00", 3071 => "00", 3072 => "00", 3073 => "00", 3074 => "00", 3075 => "00", 3076 => "00", 3077 => "00", 3078 => "00", 3079 => "00", 3080 => "00", 3081 => "00", 3082 => "00", 3083 => "00", 3084 => "00", 3085 => "00", 3086 => "00", 3087 => "00", 3088 => "00", 3089 => "00", 3090 => "00", 3091 => "00", 3092 => "00", 3093 => "00", 3094 => "00", 3095 => "00", 3096 => "00", 3097 => "00", 3098 => "00", 3099 => "00", 3100 => "00", 3101 => "00", 3102 => "00", 3103 => "00", 3104 => "00", 3105 => "00", 3106 => "00", 3107 => "00", 3108 => "00", 3109 => "00", 3110 => "00", 3111 => "00", 3112 => "00", 3113 => "00", 3114 => "00", 3115 => "00", 3116 => "00", 3117 => "00", 3118 => "00", 3119 => "00", 3120 => "00", 3121 => "00", 3122 => "00", 3123 => "00", 3124 => "00", 3125 => "00", 3126 => "00", 3127 => "00", 3128 => "00", 3129 => "00", 3130 => "00", 3131 => "00", 3132 => "00", 3133 => "00", 3134 => "00", 3135 => "00", 3136 => "00", 3137 => "00", 3138 => "00", 3139 => "00", 3140 => "00", 3141 => "00", 3142 => "00", 3143 => "00", 3144 => "00", 3145 => "00", 3146 => "00", 3147 => "00", 3148 => "00", 3149 => "00", 3150 => "00", 3151 => "00", 3152 => "00", 3153 => "00", 3154 => "00", 3155 => "00", 3156 => "00", 3157 => "00", 3158 => "00", 3159 => "00", 3160 => "00", 3161 => "00", 3162 => "00", 3163 => "00", 3164 => "00", 3165 => "00", 3166 => "00", 3167 => "00", 3168 => "00", 3169 => "00", 3170 => "00", 3171 => "00", 3172 => "00", 3173 => "00", 3174 => "00", 3175 => "00", 3176 => "00", 3177 => "00", 3178 => "00", 3179 => "00", 3180 => "00", 3181 => "00", 3182 => "00", 3183 => "00", 3184 => "00", 3185 => "00", 3186 => "00", 3187 => "00", 3188 => "00", 3189 => "00", 3190 => "00", 3191 => "00", 3192 => "00", 3193 => "00", 3194 => "00", 3195 => "00", 3196 => "00", 3197 => "00", 3198 => "00", 3199 => "00", 3200 => "00", 3201 => "00", 3202 => "00", 3203 => "00", 3204 => "00", 3205 => "00", 3206 => "00", 3207 => "00", 3208 => "00", 3209 => "00", 3210 => "00", 3211 => "00", 3212 => "00", 3213 => "00", 3214 => "00", 3215 => "00", 3216 => "00", 3217 => "00", 3218 => "00", 3219 => "00", 3220 => "00", 3221 => "00", 3222 => "00", 3223 => "00", 3224 => "00", 3225 => "00", 3226 => "00", 3227 => "00", 3228 => "00", 3229 => "00", 3230 => "00", 3231 => "00", 3232 => "00", 3233 => "00", 3234 => "00", 3235 => "00", 3236 => "00", 3237 => "00", 3238 => "00", 3239 => "00", 3240 => "00", 3241 => "00", 3242 => "00", 3243 => "00", 3244 => "00", 3245 => "00", 3246 => "00", 3247 => "00", 3248 => "00", 3249 => "00", 3250 => "00", 3251 => "00", 3252 => "00", 3253 => "00", 3254 => "00", 3255 => "00", 3256 => "00", 3257 => "00", 3258 => "00", 3259 => "00", 3260 => "00", 3261 => "00", 3262 => "00", 3263 => "00", 3264 => "00", 3265 => "00", 3266 => "00", 3267 => "00", 3268 => "00", 3269 => "00", 3270 => "00", 3271 => "00", 3272 => "00", 3273 => "00", 3274 => "00", 3275 => "00", 3276 => "00", 3277 => "00", 3278 => "00", 3279 => "00", 3280 => "00", 3281 => "00", 3282 => "00", 3283 => "00", 3284 => "00", 3285 => "00", 3286 => "00", 3287 => "00", 3288 => "00", 3289 => "00", 3290 => "00", 3291 => "00", 3292 => "00", 3293 => "00", 3294 => "00", 3295 => "00", 3296 => "00", 3297 => "00", 3298 => "00", 3299 => "00", 3300 => "00", 3301 => "00", 3302 => "00", 3303 => "00", 3304 => "00", 3305 => "00", 3306 => "00", 3307 => "00", 3308 => "00", 3309 => "00", 3310 => "00", 3311 => "00", 3312 => "00", 3313 => "00", 3314 => "00", 3315 => "00", 3316 => "00", 3317 => "00", 3318 => "00", 3319 => "00", 3320 => "00", 3321 => "00", 3322 => "00", 3323 => "00", 3324 => "00", 3325 => "00", 3326 => "00", 3327 => "00", 3328 => "00", 3329 => "00", 3330 => "00", 3331 => "00", 3332 => "00", 3333 => "00", 3334 => "00", 3335 => "00", 3336 => "00", 3337 => "00", 3338 => "00", 3339 => "00", 3340 => "00", 3341 => "00", 3342 => "00", 3343 => "00", 3344 => "00", 3345 => "00", 3346 => "00", 3347 => "00", 3348 => "00", 3349 => "00", 3350 => "00", 3351 => "00", 3352 => "00", 3353 => "00", 3354 => "00", 3355 => "00", 3356 => "00", 3357 => "00", 3358 => "00", 3359 => "00", 3360 => "00", 3361 => "00", 3362 => "00", 3363 => "00", 3364 => "00", 3365 => "00", 3366 => "00", 3367 => "00", 3368 => "00", 3369 => "00", 3370 => "00", 3371 => "00", 3372 => "00", 3373 => "00", 3374 => "00", 3375 => "00", 3376 => "00", 3377 => "00", 3378 => "00", 3379 => "00", 3380 => "00", 3381 => "00", 3382 => "00", 3383 => "00", 3384 => "00", 3385 => "00", 3386 => "00", 3387 => "00", 3388 => "00", 3389 => "00", 3390 => "00", 3391 => "00", 3392 => "00", 3393 => "00", 3394 => "00", 3395 => "00", 3396 => "00", 3397 => "00", 3398 => "00", 3399 => "00", 3400 => "00", 3401 => "00", 3402 => "00", 3403 => "00", 3404 => "00", 3405 => "00", 3406 => "00", 3407 => "00", 3408 => "00", 3409 => "00", 3410 => "00", 3411 => "00", 3412 => "00", 3413 => "00", 3414 => "00", 3415 => "00", 3416 => "00", 3417 => "00", 3418 => "00", 3419 => "00", 3420 => "00", 3421 => "00", 3422 => "00", 3423 => "00", 3424 => "00", 3425 => "00", 3426 => "00", 3427 => "00", 3428 => "00", 3429 => "00", 3430 => "00", 3431 => "00", 3432 => "00", 3433 => "00", 3434 => "00", 3435 => "00", 3436 => "00", 3437 => "00", 3438 => "00", 3439 => "00", 3440 => "00", 3441 => "00", 3442 => "00", 3443 => "00", 3444 => "00", 3445 => "00", 3446 => "00", 3447 => "00", 3448 => "00", 3449 => "00", 3450 => "00", 3451 => "00", 3452 => "00", 3453 => "00", 3454 => "00", 3455 => "00", 3456 => "00", 3457 => "00", 3458 => "00", 3459 => "00", 3460 => "00", 3461 => "00", 3462 => "00", 3463 => "00", 3464 => "00", 3465 => "00", 3466 => "00", 3467 => "00", 3468 => "00", 3469 => "00", 3470 => "00", 3471 => "00", 3472 => "00", 3473 => "00", 3474 => "00", 3475 => "00", 3476 => "00", 3477 => "00", 3478 => "00", 3479 => "00", 3480 => "00", 3481 => "00", 3482 => "00", 3483 => "00", 3484 => "00", 3485 => "00", 3486 => "00", 3487 => "00", 3488 => "00", 3489 => "00", 3490 => "00", 3491 => "00", 3492 => "00", 3493 => "00", 3494 => "00", 3495 => "00", 3496 => "00", 3497 => "00", 3498 => "00", 3499 => "00", 3500 => "00", 3501 => "00", 3502 => "00", 3503 => "00", 3504 => "00", 3505 => "00", 3506 => "00", 3507 => "00", 3508 => "00", 3509 => "00", 3510 => "00", 3511 => "00", 3512 => "00", 3513 => "00", 3514 => "00", 3515 => "00", 3516 => "00", 3517 => "00", 3518 => "00", 3519 => "00", 3520 => "00", 3521 => "00", 3522 => "00", 3523 => "00", 3524 => "00", 3525 => "00", 3526 => "00", 3527 => "00", 3528 => "00", 3529 => "00", 3530 => "00", 3531 => "00", 3532 => "00", 3533 => "00", 3534 => "00", 3535 => "00", 3536 => "00", 3537 => "00", 3538 => "00", 3539 => "00", 3540 => "00", 3541 => "00", 3542 => "00", 3543 => "00", 3544 => "00", 3545 => "00", 3546 => "00", 3547 => "00", 3548 => "00", 3549 => "00", 3550 => "00", 3551 => "00", 3552 => "00", 3553 => "00", 3554 => "00", 3555 => "00", 3556 => "00", 3557 => "00", 3558 => "00", 3559 => "00", 3560 => "00", 3561 => "00", 3562 => "00", 3563 => "00", 3564 => "00", 3565 => "00", 3566 => "00", 3567 => "00", 3568 => "00", 3569 => "00", 3570 => "00", 3571 => "00", 3572 => "00", 3573 => "00", 3574 => "00", 3575 => "00", 3576 => "00", 3577 => "00", 3578 => "00", 3579 => "00", 3580 => "00", 3581 => "00", 3582 => "00", 3583 => "00", 3584 => "00", 3585 => "00", 3586 => "00", 3587 => "00", 3588 => "00", 3589 => "00", 3590 => "00", 3591 => "00", 3592 => "00", 3593 => "00", 3594 => "00", 3595 => "00", 3596 => "00", 3597 => "00", 3598 => "00", 3599 => "00", 3600 => "00", 3601 => "00", 3602 => "00", 3603 => "00", 3604 => "00", 3605 => "00", 3606 => "00", 3607 => "00", 3608 => "00", 3609 => "00", 3610 => "00", 3611 => "00", 3612 => "00", 3613 => "00", 3614 => "00", 3615 => "00", 3616 => "00", 3617 => "00", 3618 => "00", 3619 => "00", 3620 => "00", 3621 => "00", 3622 => "00", 3623 => "00", 3624 => "00", 3625 => "00", 3626 => "00", 3627 => "00", 3628 => "00", 3629 => "00", 3630 => "00", 3631 => "00", 3632 => "00", 3633 => "00", 3634 => "00", 3635 => "00", 3636 => "00", 3637 => "00", 3638 => "00", 3639 => "00", 3640 => "00", 3641 => "00", 3642 => "00", 3643 => "00", 3644 => "00", 3645 => "00", 3646 => "00", 3647 => "00", 3648 => "00", 3649 => "00", 3650 => "00", 3651 => "00", 3652 => "00", 3653 => "00", 3654 => "00", 3655 => "00", 3656 => "00", 3657 => "00", 3658 => "00", 3659 => "00", 3660 => "00", 3661 => "00", 3662 => "00", 3663 => "00", 3664 => "00", 3665 => "00", 3666 => "00", 3667 => "00", 3668 => "00", 3669 => "00", 3670 => "00", 3671 => "00", 3672 => "00", 3673 => "00", 3674 => "00", 3675 => "00", 3676 => "00", 3677 => "00", 3678 => "00", 3679 => "00", 3680 => "00", 3681 => "00", 3682 => "00", 3683 => "00", 3684 => "00", 3685 => "00", 3686 => "00", 3687 => "00", 3688 => "00", 3689 => "00", 3690 => "00", 3691 => "00", 3692 => "00", 3693 => "00", 3694 => "00", 3695 => "00", 3696 => "00", 3697 => "00", 3698 => "00", 3699 => "00", 3700 => "00", 3701 => "00", 3702 => "00", 3703 => "00", 3704 => "00", 3705 => "00", 3706 => "00", 3707 => "00", 3708 => "00", 3709 => "00", 3710 => "00", 3711 => "00", 3712 => "00", 3713 => "00", 3714 => "00", 3715 => "00", 3716 => "00", 3717 => "00", 3718 => "00", 3719 => "00", 3720 => "00", 3721 => "00", 3722 => "00", 3723 => "00", 3724 => "00", 3725 => "00", 3726 => "00", 3727 => "00", 3728 => "00", 3729 => "00", 3730 => "00", 3731 => "00", 3732 => "00", 3733 => "00", 3734 => "00", 3735 => "00", 3736 => "00", 3737 => "00", 3738 => "00", 3739 => "00", 3740 => "00", 3741 => "00", 3742 => "00", 3743 => "00", 3744 => "00", 3745 => "00", 3746 => "00", 3747 => "00", 3748 => "00", 3749 => "00", 3750 => "00", 3751 => "00", 3752 => "00", 3753 => "00", 3754 => "00", 3755 => "00", 3756 => "00", 3757 => "00", 3758 => "00", 3759 => "00", 3760 => "00", 3761 => "00", 3762 => "00", 3763 => "00", 3764 => "00", 3765 => "00", 3766 => "00", 3767 => "00", 3768 => "00", 3769 => "00", 3770 => "00", 3771 => "00", 3772 => "00", 3773 => "00", 3774 => "01", 3775 => "11", 3776 => "10", 3777 => "11", 3778 => "01", 3779 => "11", 3780 => "01", 3781 => "00", 3782 => "10", 3783 => "11", 3784 => "10", 3785 => "11", 3786 => "01", 3787 => "11", 3788 => "01", 3789 => "00", 3790 => "10", 3791 => "11", 3792 => "10", 3793 => "11", 3794 => "01", 3795 => "11", 3796 => "01", 3797 => "00", 3798 => "10", 3799 => "11", 3800 => "01", 3801 => "00", 3802 => "10", 3803 => "00", 3804 => "01", 3805 => "11", 3806 => "01", 3807 => "11", 3808 => "01", 3809 => "11", 3810 => "10", 3811 => "11", 3812 => "01", 3813 => "00", 3814 => "01", 3815 => "11", 3816 => "10", 3817 => "00", 3818 => "10", 3819 => "11", 3820 => "10", 3821 => "11", 3822 => "10", 3823 => "00", 3824 => "01", 3825 => "11", 3826 => "10", 3827 => "11", 3828 => "01", 3829 => "00", 3830 => "10", 3831 => "00", 3832 => "10", 3833 => "00", 3834 => "01", 3835 => "11", 3836 => "10", 3837 => "00", 3838 => "10", 3839 => "11", 3840 => "01", 3841 => "00", 3842 => "10", 3843 => "00", 3844 => "01", 3845 => "11", 3846 => "10", 3847 => "00", 3848 => "01", 3849 => "11", 3850 => "01", 3851 => "00", 3852 => "10", 3853 => "11", 3854 => "01", 3855 => "11", others => "00");
	
	-- Adresse som peger på den ROM-plads der skal læses fra
    signal address : integer range 0 to ROM_SIZE - 1 := 0;

begin

    -- Main process: Læser ROM-værdi ved rising_edge af clk og outputter dette som data og strobe
    process(clk50mhz )
    begin
        if rising_edge(clk50mhz ) then
            if reset = '1' then
                address     <= 0;
                D    <= '0';
                S    <= '0';
            else
                D    <= rom(address)(1);
                S    <= rom(address)(0);
                address     <= address + 1;
            end if;
        end if;
    end process;

end architecture;
